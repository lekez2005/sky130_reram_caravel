// Generated from OpenRAM

module reram_sram1 (
    INPUT [6:0] addr,
    INPUT clk,
    INPUT csb,
    INPUT [6:0] data,
    INPUT data_others,
    OUTPUT [6:0] data_out,
    INOUT gnd,
    INPUT [6:0] mask,
    INPUT mask_others,
    INPUT sense_trig,
    INPUT vclamp,
    INPUT vclampp,
    INOUT vdd,
    INOUT vdd_wordline,
    INOUT vdd_write,
    INPUT vref,
    INPUT web,
);
