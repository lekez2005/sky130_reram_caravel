.subckt sky130_fd_pr__reram_reram_cell TE BE
.ends
